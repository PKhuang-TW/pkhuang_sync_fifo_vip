`ifndef FIFO_DEFINE_SVH
`define FIFO_DEFINE_SVH

`define     D_DATA_WIDTH    8
`define     D_FIFO_DEPTH    16
`define     D_ADDR_WIDTH    $clog2(`D_FIFO_DEPTH)

`endif