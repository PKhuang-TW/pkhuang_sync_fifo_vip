`ifndef FIFO_DEFINE_SVH
`define FIFO_DEFINE_SVH

parameter   P_DATA_WIDTH  = 8;
parameter   P_FIFO_DEPTH  = 16;

`endif