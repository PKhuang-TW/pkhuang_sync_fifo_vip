`ifndef FIFO_PACKAGE_SVH
`define FIFO_PACKAGE_SVH

package fifo_package;
    parameter   P_DATA_WIDTH  = 8;
    parameter   P_FIFO_DEPTH  = 16;
endpackage

`endif